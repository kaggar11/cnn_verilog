`timescale 1ns/1ps
module InputPad_tb;

// Inputs
       
  		parameter SIZE=7;
  		parameter FILTER_SIZE=3;
  		parameter size=SIZE;
  		parameter filter_size=FILTER_SIZE;
 // logic [31:0] outputsize1;
  //parameter outputsize= SIZE+FILTER_SIZE-(SIZE%FILTER_SIZE);
 // parameter outputsize= SIZE-((SIZE%FILTER_SIZE)-(FILTER_SIZE));
  parameter outputsize=SIZE+(((FILTER_SIZE-(SIZE%FILTER_SIZE)))%FILTER_SIZE);
  //arameter outputsize=SIZE+FILTER_SIZE-(SIZE%FILTER_SIZE);
  logic [31:0] array1[0:(SIZE-1)][0:(SIZE-1)];
  logic [31:0] array2[0:(outputsize-1)][0:(outputsize-1)];
  logic clk;
  logic en;
  logic reset;
  //parameter outputsize=(2*(size-1))+1;
// Outputs
  int row;
  int col;
// Instantiate the Unit Under Test (UUT)
  InputPad #(.SIZE(size),.FILTER_SIZE(filter_size)) uut(.clk(clk),.en(en),.reset(reset),.array1(array1),.array2(array2));
  


  
  
		initial begin
// Initialize Inputs
          $display("Starting ghfhgfhgfh");
          //$display("This is outputsize:%0d",outputsize);
          //$finish;
			clk = 0;
			en = 0;
			reset = 1;
              for(row=0;row<size;row=row+1) begin 
                for(col=0;col<size;col=col+1) begin 
                  array1[row][col]='d3;
                  $display("array1[%d][%d]=%0d", row,col,array1[row][col]);
      			    end 
    		    end
          $display("Hellrtetretertreo");
            @(posedge clk);
             reset=0;
             en=1;
          @(posedge clk);
          $display("gfgfgf");
           #9000
          for(row=0;row<outputsize;row=row+1) begin 
            for(col=0;col<outputsize;col=col+1)  begin 
             // $display("This is row=%0d and col=%0d",row,col);
              $display("This is array2[%0d][%0d]=%0d",row,col,array2[row][col]);
            end 
          end 
          //  $finish;
         ;
          $finish;
           end
  
  
//blocks_in[0+:4][0+:3][0+:3] = 0;

// Wait 100 ns for global reset to finish
//#5000;
//       end
// Add stimulus here
           always begin
			#250 clk=!clk;
			end
//initial begin
//@(posedge clk);
//control=1;
//reset  =0;
//blocks_in[0][0+:3][0+:3] = 64'b1;
//end
     
endmodule
